// +FHDR============================================================================/
// Author       : mayia
// Creat Time   : 2020/07/14 11:47:10
// File Name    : inst_tx_top.v
// Module Ver   : Vx.x
//
//
// All Rights Reserved
//
// ---------------------------------------------------------------------------------/
//
// Modification History:
// V1.0         initial
//
// -FHDR============================================================================/
// 
// inst_tx_ctrl
//    |---
// 
`timescale 1ns/1ps

module inst_tx_top #
(
    parameter                       U_DLY = 1                   
)
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    input                           clk_sys                     , 
    input                           rst_n                       , 
// ----------------------------------------------------------------------------
// Config Register Data
// ----------------------------------------------------------------------------
    input                    [15:0] cfg_ins_txcnt               , // 指令发送次数
    input                    [15:0] cfg_ins_length              , // 指令长度
    input                    [31:0] cfg_ins_waittime            , // 发送间隔时间
    input                           cfg_keyer_sel               , // 调制体制选择  
// ----------------------------------------------------------------------------
// Time
// ----------------------------------------------------------------------------
    input                    [63:0] local_time                  , 
// ----------------------------------------------------------------------------
// Instruct Data From Memory
// ----------------------------------------------------------------------------
    input                   [511:0] inst_data                   , 
    input                           inst_data_valid             , 
// ----------------------------------------------------------------------------
// Log Instruct Data 
// ----------------------------------------------------------------------------
    output                  [575:0] log_inst_data               , 
    output                          log_inst_data_valid         , 
// ----------------------------------------------------------------------------
// PCM Instruct Data
// ----------------------------------------------------------------------------
    output                  [511:0] pcm_tx_data                 , 
    output                          pcm_tx_data_valid           , 
// ----------------------------------------------------------------------------
// DY Instruct Data
// ----------------------------------------------------------------------------
    output                  [127:0] dy_tx_data                  , 
    output                          dy_tx_data_valid            , 
// ----------------------------------------------------------------------------
// Debug Status
// ----------------------------------------------------------------------------
    output                          debug_tx_overflow             
);

wire                        [511:0] pcm_inst_data               ; 
wire                                pcm_inst_data_valid         ; 

wire                        [511:0] dy_inst_data                ; 
wire                                dy_inst_data_valid          ; 

inst_tx_ctrl #
(
    .U_DLY                          (U_DLY                      )  
)
u_inst_tx_ctrl
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Config Register Data
// ----------------------------------------------------------------------------
    .cfg_ins_txcnt                  (cfg_ins_txcnt[15:0]        ), // (input ) 指令发送次数
    .cfg_ins_waittime               (cfg_ins_waittime[31:0]     ), // (input ) 发送间隔时间
    .cfg_keyer_sel                  (cfg_keyer_sel              ), // (input )调制体制选择  
// ----------------------------------------------------------------------------
// Time
// ----------------------------------------------------------------------------
    .local_time                     (local_time[63:0]           ), // (input )
// ----------------------------------------------------------------------------
// Instruct Data From Memory
// ----------------------------------------------------------------------------
    .inst_data                      (inst_data[511:0]           ), // (input )
    .inst_data_valid                (inst_data_valid            ), // (input )
// ----------------------------------------------------------------------------
// Log TX Data
// ----------------------------------------------------------------------------
    .log_inst_data                  (log_inst_data[575:0]       ), // (output)
    .log_inst_data_valid            (log_inst_data_valid        ), // (output)
// ----------------------------------------------------------------------------
// PCM TX Data
// ----------------------------------------------------------------------------
    .pcm_inst_data                  (pcm_inst_data[511:0]       ), // (output)
    .pcm_inst_data_valid            (pcm_inst_data_valid        ), // (output)
// ----------------------------------------------------------------------------
// DY TX Data
// ----------------------------------------------------------------------------
    .dy_inst_data                   (dy_inst_data[511:0]        ), // (output)
    .dy_inst_data_valid             (dy_inst_data_valid         ), // (output)
// ----------------------------------------------------------------------------
// Debug Status
// ----------------------------------------------------------------------------
    .debug_tx_overflow              (debug_tx_overflow          )  // (output)
);

inst_tx2pcm #
(
    .U_DLY                          (U_DLY                      )  
)
u_inst_tx2pcm
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Config Register Data
// ----------------------------------------------------------------------------
    .cfg_ins_length                 (cfg_ins_length[15:0]       ), // (input ) 指令长度
// ----------------------------------------------------------------------------
// PCM TX Control
// ----------------------------------------------------------------------------
    .pcm_inst_data                  (pcm_inst_data[511:0]       ), // (input )
    .pcm_inst_data_valid            (pcm_inst_data_valid        ), // (input )
// ----------------------------------------------------------------------------
// PCM Instruct Data
// ----------------------------------------------------------------------------
    .pcm_tx_data                    (pcm_tx_data[511:0]         ), // (output)
    .pcm_tx_data_valid              (pcm_tx_data_valid          )  // (output)
);

inst_tx2dy #
(
    .U_DLY                          (U_DLY                      )  
)
u_inst_tx2dy
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Config Register Data
// ----------------------------------------------------------------------------
    .cfg_ins_length                 (cfg_ins_length[15:0]       ), // (input ) 指令长度
// ----------------------------------------------------------------------------
// PCM TX Control
// ----------------------------------------------------------------------------
    .dy_inst_data                   (dy_inst_data[511:0]        ), // (input )
    .dy_inst_data_valid             (dy_inst_data_valid         ), // (input )
// ----------------------------------------------------------------------------
// PCM Instruct Data
// ----------------------------------------------------------------------------
    .dy_tx_data                     (dy_tx_data[127:0]          ), // (output)
    .dy_tx_data_valid               (dy_tx_data_valid           )  // (output)
);

endmodule



