// +FHDR============================================================================/
// Author       : mayia
// Creat Time   : 2020/07/14 17:28:18
// File Name    : key_top.v
// Module Ver   : Vx.x
//
//
// All Rights Reserved
//
// ---------------------------------------------------------------------------------/
//
// Modification History:
// V1.0         initial
//
// -FHDR============================================================================/
// 
// key_top
//    |---
// 
`timescale 1ns/1ps

module key_top #
(
    parameter                       U_DLY = 1
)
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    input                           clk_sys                     , 
    input                           rst_n                       , 
// ----------------------------------------------------------------------------
// Config
// ----------------------------------------------------------------------------
    input                    [31:0] cfg_key_filter_data         , 
// ----------------------------------------------------------------------------
// Key In
// ----------------------------------------------------------------------------
    input                    [15:0] key_in                      , 
// ----------------------------------------------------------------------------
// Key Data
// ----------------------------------------------------------------------------
    output                   [15:0] key_data                    , 
    output                          key_data_valid              ,

    output                          key_lr_status               , 
    output                          key_status_valid            , 
// ----------------------------------------------------------------------------
// Key Instruct
// ----------------------------------------------------------------------------
    output                          key_instruct_valid          , 
    output                   [15:0] key_instruct                  
);

wire                         [15:0] key_edge_r                  ; 
wire                         [15:0] key_edge_f                  ; 
wire                         [15:0] key_edge_rf                 ; 

genvar                              i,j                         ;

generate
for(i=0;i<16;i=i+1)
begin:filter_loop
cb_line_filter #
(
    .U_DLY                          (U_DLY                      )  
)
u_cb_line_filter
( 
//-----------------------------------------------------------------------------------
// Golbal Signals
//-----------------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
//-----------------------------------------------------------------------------------
// filter paramter
//-----------------------------------------------------------------------------------
    .filter_cnt                     (cfg_key_filter_data[31:0]  ), // (input ) 
//-----------------------------------------------------------------------------------
// line signal
//-----------------------------------------------------------------------------------
    .sig_in                         (key_in[i]                  ), // (input )
    .sig_out                        (key_data[i]                )  // (output)
);
end
endgenerate

generate
for(j=0;j<16;j=j+1)
begin:edge_loop
cb_edge_cap #
(
    .U_DLY                          (U_DLY                      )  
)
u_cb_edge_cap
(
//-----------------------------------------------------------------------------------
// Golbal Signals
//-----------------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
//-----------------------------------------------------------------------------------
// signal in
//-----------------------------------------------------------------------------------
    .sig_in                         (key_data[j]                ), // (input )
//-----------------------------------------------------------------------------------
// Result Signals
//-----------------------------------------------------------------------------------
    .edge_r                         (key_edge_r[j]              ), // (output)
    .edge_f                         (key_edge_f[j]              ), // (output)
    .edge_rf                        (key_edge_rf[j]             )  // (output)
);
end
endgenerate

assign key_data_valid = |key_edge_f[4:0];
assign key_status_valid = key_edge_rf[5];
assign key_lr_status = key_data[5];

key_deframe #
(
    .U_DLY                          (U_DLY                      )  
)
u_key_deframe
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Key Data
// ----------------------------------------------------------------------------
    .key_data                       (key_data[15:0]             ), // (input )
    .key_data_valid                 (key_data_valid             ), // (input )
// ----------------------------------------------------------------------------
// Key Instruct
// ----------------------------------------------------------------------------
    .key_instruct                   (key_instruct[15:0]         ), // (output)
    .key_instruct_valid             (key_instruct_valid         )  // (output)
);

endmodule



