// +FHDR============================================================================/
// Author       : mayia
// Creat Time   : 2020/07/14 10:17:39
// File Name    : uart_top.v
// Module Ver   : Vx.x
//
//
// All Rights Reserved
//
// ---------------------------------------------------------------------------------/
//
// Modification History:
// V1.0         initial
//
// -FHDR============================================================================/
// 
// uart_top
//    |---
// 
`timescale 1ns/1ps

module uart_top #
(
    parameter                       U_DLY = 1
)
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    input                           clk_sys                     , 
    input                           rst_n                       , 
//-----------------------------------------------------------------------------
// Config Port
//-----------------------------------------------------------------------------
    input                    [15:0] baud_rate                   , 
    input                     [3:0] data_width                  , 
    input                           check_en                    , 
    input                           check_sel                   , 
    input                           check_filter                , 
    input                           stop_bit                    , 
// ----------------------------------------------------------------------------
// Send Data 
// ----------------------------------------------------------------------------
    input                           uart_tx_en                  , 
    input                     [7:0] uart_tx_data                , 
// ----------------------------------------------------------------------------
// Receive Data
// ----------------------------------------------------------------------------
    output                    [7:0] uart_rx_data                , 
    output                          uart_rx_data_valid          , 
// ----------------------------------------------------------------------------
// Uart
// ----------------------------------------------------------------------------
    input                           uart_rx                     , 
    output                          uart_tx                       
);

wire                                baud_en                     ; 

wire                                fifo_rd_en                  ; 
wire                          [7:0] fifo_rd_data                ; 
wire                                fifo_empty                  ; 

wire                                tx_busy                     ; 

wire                          [7:0] driver_tx_data              ; 
wire                                driver_tx_data_valid        ; 

uart_baud #
(
    .U_DLY                          (U_DLY                      ), 
    .DW                             (16                         )  
)
u_uart_baud
(
//-----------------------------------------------------------------------------------
// Clock & Reset
//-----------------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
//-----------------------------------------------------------------------------------
// Other Signals
//-----------------------------------------------------------------------------------
    .baud_rate                      (baud_rate[15:0]            ), // (input )
    .baud_en                        (baud_en                    )  // (output)
);

fifo_d1kw8_st	u_fifo_d1kw8_st
(
    .aclr                           (!rst_n                     ), 
    .clock                          (clk_sys                    ), 
    .wrreq                          (uart_tx_en                 ), 
    .data                           (uart_tx_data[7:0]          ), 
    .rdreq                          (fifo_rd_en                 ), 
    .q                              (fifo_rd_data[7:0]          ), 
    .empty                          (fifo_empty                 ), 
    .full                           (                           ), 
    .usedw                          (/* not used */             )  
);

uart_txctrl #
(
    .U_DLY                          (U_DLY                      )  
)
u_uart_txctrl
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// FIFO Read 
// ----------------------------------------------------------------------------
    .fifo_rd_en                     (fifo_rd_en                 ), // (output)
    .fifo_rd_data                   (fifo_rd_data[7:0]          ), // (input )
    .fifo_empty                     (fifo_empty                 ), // (input )
// ----------------------------------------------------------------------------
// Send status
// ----------------------------------------------------------------------------
    .tx_busy                        (tx_busy                    ), // (input )
// ----------------------------------------------------------------------------
// Send Data 
// ----------------------------------------------------------------------------
    .driver_tx_data                 (driver_tx_data[7:0]        ), // (output)
    .driver_tx_data_valid           (driver_tx_data_valid       )  // (output)
);

uart_tx #
(
    .U_DLY                          (U_DLY                      )  
)
u_uart_tx
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Config Data 
// ----------------------------------------------------------------------------
    .baud_en                        (baud_en                    ), // (input )

    .data_width                     (data_width[3:0]            ), // (input )
    .check_en                       (check_en                   ), // (input )
    .check_sel                      (check_sel                  ), // (input )
    .stop_bit                       (stop_bit                   ), // (input )

    .tx_busy                        (tx_busy                    ), // (output)
// ----------------------------------------------------------------------------
// Send Data 
// ----------------------------------------------------------------------------
    .driver_tx_data                 (driver_tx_data[7:0]        ), // (input )
    .driver_tx_data_valid           (driver_tx_data_valid       ), // (input )
// ----------------------------------------------------------------------------
// Uart
// ----------------------------------------------------------------------------
    .uart_tx                        (uart_tx                    )  // (output)
);

uart_rx #
(
    .U_DLY                          (U_DLY                      )  
)
u_uart_rx
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Config Data 
// ----------------------------------------------------------------------------
    .baud_en                        (baud_en                    ), // (input )

    .data_width                     (data_width[3:0]            ), // (input )
    .check_en                       (check_en                   ), // (input )
    .check_sel                      (check_sel                  ), // (input )
    .check_filter                   (check_filter               ), // (input )
    .stop_bit                       (stop_bit                   ), // (input )
// ----------------------------------------------------------------------------
// Uart
// ----------------------------------------------------------------------------
    .uart_rx                        (uart_rx                    ), // (input )
// ----------------------------------------------------------------------------
// Receive Data 
// ----------------------------------------------------------------------------
    .driver_rx_data                 (uart_rx_data[7:0]          ), // (output)
    .driver_rx_data_valid           (uart_rx_data_valid         ), // (output)
// ----------------------------------------------------------------------------
// Debug
// ----------------------------------------------------------------------------
    .debug_check_error              (                           ), // (output)
    .debug_stop_error               (                           )  // (output)
);

endmodule




