// +FHDR============================================================================/
// Author       : huangjie
// Creat Time   : 2020/08/05 18:48:21
// File Name    : dymodem_test.v
// Module Ver   : Vx.x
//
//
// All Rights Reserved
//
// ---------------------------------------------------------------------------------/
//
// Modification History:
// V1.0         initial
//
// -FHDR============================================================================/
// 
// dymodem_test
//    |---
// 
`timescale 1ns/1ps

module dymodem_test ;


reg                                 clk_sys                     ; 
reg                                 rst_n                       ; 

wire                        [127:0] dy_tx_data                  ; 

assign dy_tx_data = 128'h0001_1e00_01e0_001e_1e00_01e0_001e_1e00;

wire                         [11:0] dy_idata                    ; 
wire                         [11:0] dy_qdata                    ; 

iqmodem_dy #
(
    .U_DLY                          (1                          )  
)
u_iqmodem_dy
(
// ----------------------------------------------------------------------------
// Clock & Reset
// ----------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ----------------------------------------------------------------------------
// Config
// ----------------------------------------------------------------------------
    .cfg_dy_load_en                 (1'b1                       ), // (input )
    .cfg_dy_keyer_en                (1'b1                       ), // (input )
    .cfg_dy_fbias                   (16'd50                     ), // (input )
// ----------------------------------------------------------------------------
// DY Instruct Data
// ----------------------------------------------------------------------------
    .dy_tx_en                       (1'b1                       ), // (input )
    .dy_tx_data                     (dy_tx_data[127:0]          ), // (input )
// ----------------------------------------------------------------------------
// DAC data
// ----------------------------------------------------------------------------
    .dy_idata                       (dy_idata[11:0]             ), // (output)
    .dy_qdata                       (dy_qdata[11:0]             )  // (output)
);


initial 
begin
    clk_sys = 0;
    rst_n = 0;

    #100;
    rst_n = 1;
end

always #8  clk_sys = ~clk_sys;

endmodule   





